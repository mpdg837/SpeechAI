module hamming_window_array(
	input clk,
	input rst,
	
	input[8:0] mul_addr,
	output reg[15:0] mul_out
);


reg[15:0] multiplies[511:0];
initial begin
	multiplies[0]=5027;
	multiplies[1]=5030;
	multiplies[2]=5036;
	multiplies[3]=5048;
	multiplies[4]=5064;
	multiplies[5]=5085;
	multiplies[6]=5110;
	multiplies[7]=5139;
	multiplies[8]=5174;
	multiplies[9]=5212;
	multiplies[10]=5256;
	multiplies[11]=5304;
	multiplies[12]=5356;
	multiplies[13]=5413;
	multiplies[14]=5474;
	multiplies[15]=5540;
	multiplies[16]=5611;
	multiplies[17]=5686;
	multiplies[18]=5765;
	multiplies[19]=5849;
	multiplies[20]=5938;
	multiplies[21]=6030;
	multiplies[22]=6128;
	multiplies[23]=6229;
	multiplies[24]=6335;
	multiplies[25]=6445;
	multiplies[26]=6560;
	multiplies[27]=6679;
	multiplies[28]=6803;
	multiplies[29]=6930;
	multiplies[30]=7062;
	multiplies[31]=7199;
	multiplies[32]=7339;
	multiplies[33]=7484;
	multiplies[34]=7633;
	multiplies[35]=7786;
	multiplies[36]=7943;
	multiplies[37]=8105;
	multiplies[38]=8270;
	multiplies[39]=8440;
	multiplies[40]=8613;
	multiplies[41]=8791;
	multiplies[42]=8973;
	multiplies[43]=9158;
	multiplies[44]=9348;
	multiplies[45]=9542;
	multiplies[46]=9739;
	multiplies[47]=9940;
	multiplies[48]=10145;
	multiplies[49]=10354;
	multiplies[50]=10567;
	multiplies[51]=10783;
	multiplies[52]=11004;
	multiplies[53]=11227;
	multiplies[54]=11455;
	multiplies[55]=11686;
	multiplies[56]=11920;
	multiplies[57]=12159;
	multiplies[58]=12400;
	multiplies[59]=12645;
	multiplies[60]=12894;
	multiplies[61]=13146;
	multiplies[62]=13401;
	multiplies[63]=13659;
	multiplies[64]=13921;
	multiplies[65]=14186;
	multiplies[66]=14455;
	multiplies[67]=14726;
	multiplies[68]=15000;
	multiplies[69]=15278;
	multiplies[70]=15559;
	multiplies[71]=15842;
	multiplies[72]=16129;
	multiplies[73]=16418;
	multiplies[74]=16710;
	multiplies[75]=17005;
	multiplies[76]=17303;
	multiplies[77]=17604;
	multiplies[78]=17907;
	multiplies[79]=18213;
	multiplies[80]=18521;
	multiplies[81]=18832;
	multiplies[82]=19146;
	multiplies[83]=19462;
	multiplies[84]=19780;
	multiplies[85]=20100;
	multiplies[86]=20423;
	multiplies[87]=20749;
	multiplies[88]=21076;
	multiplies[89]=21405;
	multiplies[90]=21737;
	multiplies[91]=22071;
	multiplies[92]=22406;
	multiplies[93]=22744;
	multiplies[94]=23083;
	multiplies[95]=23425;
	multiplies[96]=23768;
	multiplies[97]=24113;
	multiplies[98]=24459;
	multiplies[99]=24807;
	multiplies[100]=25157;
	multiplies[101]=25509;
	multiplies[102]=25861;
	multiplies[103]=26216;
	multiplies[104]=26571;
	multiplies[105]=26928;
	multiplies[106]=27286;
	multiplies[107]=27646;
	multiplies[108]=28006;
	multiplies[109]=28368;
	multiplies[110]=28730;
	multiplies[111]=29094;
	multiplies[112]=29459;
	multiplies[113]=29824;
	multiplies[114]=30190;
	multiplies[115]=30557;
	multiplies[116]=30925;
	multiplies[117]=31294;
	multiplies[118]=31663;
	multiplies[119]=32032;
	multiplies[120]=32402;
	multiplies[121]=32773;
	multiplies[122]=33144;
	multiplies[123]=33515;
	multiplies[124]=33886;
	multiplies[125]=34258;
	multiplies[126]=34630;
	multiplies[127]=35002;
	multiplies[128]=35374;
	multiplies[129]=35746;
	multiplies[130]=36118;
	multiplies[131]=36490;
	multiplies[132]=36861;
	multiplies[133]=37233;
	multiplies[134]=37604;
	multiplies[135]=37974;
	multiplies[136]=38345;
	multiplies[137]=38714;
	multiplies[138]=39084;
	multiplies[139]=39453;
	multiplies[140]=39821;
	multiplies[141]=40188;
	multiplies[142]=40555;
	multiplies[143]=40921;
	multiplies[144]=41286;
	multiplies[145]=41650;
	multiplies[146]=42013;
	multiplies[147]=42375;
	multiplies[148]=42736;
	multiplies[149]=43096;
	multiplies[150]=43455;
	multiplies[151]=43812;
	multiplies[152]=44169;
	multiplies[153]=44524;
	multiplies[154]=44877;
	multiplies[155]=45229;
	multiplies[156]=45580;
	multiplies[157]=45929;
	multiplies[158]=46276;
	multiplies[159]=46622;
	multiplies[160]=46966;
	multiplies[161]=47308;
	multiplies[162]=47648;
	multiplies[163]=47987;
	multiplies[164]=48324;
	multiplies[165]=48658;
	multiplies[166]=48991;
	multiplies[167]=49321;
	multiplies[168]=49650;
	multiplies[169]=49976;
	multiplies[170]=50300;
	multiplies[171]=50622;
	multiplies[172]=50941;
	multiplies[173]=51259;
	multiplies[174]=51573;
	multiplies[175]=51885;
	multiplies[176]=52195;
	multiplies[177]=52502;
	multiplies[178]=52807;
	multiplies[179]=53109;
	multiplies[180]=53408;
	multiplies[181]=53704;
	multiplies[182]=53998;
	multiplies[183]=54289;
	multiplies[184]=54577;
	multiplies[185]=54862;
	multiplies[186]=55144;
	multiplies[187]=55423;
	multiplies[188]=55699;
	multiplies[189]=55972;
	multiplies[190]=56242;
	multiplies[191]=56508;
	multiplies[192]=56772;
	multiplies[193]=57032;
	multiplies[194]=57289;
	multiplies[195]=57543;
	multiplies[196]=57793;
	multiplies[197]=58040;
	multiplies[198]=58283;
	multiplies[199]=58523;
	multiplies[200]=58759;
	multiplies[201]=58992;
	multiplies[202]=59221;
	multiplies[203]=59447;
	multiplies[204]=59669;
	multiplies[205]=59887;
	multiplies[206]=60102;
	multiplies[207]=60312;
	multiplies[208]=60519;
	multiplies[209]=60723;
	multiplies[210]=60922;
	multiplies[211]=61118;
	multiplies[212]=61309;
	multiplies[213]=61497;
	multiplies[214]=61680;
	multiplies[215]=61860;
	multiplies[216]=62036;
	multiplies[217]=62207;
	multiplies[218]=62375;
	multiplies[219]=62538;
	multiplies[220]=62698;
	multiplies[221]=62853;
	multiplies[222]=63004;
	multiplies[223]=63151;
	multiplies[224]=63293;
	multiplies[225]=63432;
	multiplies[226]=63566;
	multiplies[227]=63696;
	multiplies[228]=63821;
	multiplies[229]=63943;
	multiplies[230]=64060;
	multiplies[231]=64172;
	multiplies[232]=64280;
	multiplies[233]=64384;
	multiplies[234]=64483;
	multiplies[235]=64578;
	multiplies[236]=64669;
	multiplies[237]=64755;
	multiplies[238]=64837;
	multiplies[239]=64914;
	multiplies[240]=64987;
	multiplies[241]=65055;
	multiplies[242]=65119;
	multiplies[243]=65178;
	multiplies[244]=65233;
	multiplies[245]=65283;
	multiplies[246]=65328;
	multiplies[247]=65369;
	multiplies[248]=65406;
	multiplies[249]=65438;
	multiplies[250]=65465;
	multiplies[251]=65488;
	multiplies[252]=65506;
	multiplies[253]=65520;
	multiplies[254]=65529;
	multiplies[255]=65534;
	multiplies[256]=65534;
	multiplies[257]=65529;
	multiplies[258]=65520;
	multiplies[259]=65506;
	multiplies[260]=65488;
	multiplies[261]=65465;
	multiplies[262]=65438;
	multiplies[263]=65406;
	multiplies[264]=65369;
	multiplies[265]=65328;
	multiplies[266]=65283;
	multiplies[267]=65233;
	multiplies[268]=65178;
	multiplies[269]=65119;
	multiplies[270]=65055;
	multiplies[271]=64987;
	multiplies[272]=64914;
	multiplies[273]=64837;
	multiplies[274]=64755;
	multiplies[275]=64669;
	multiplies[276]=64578;
	multiplies[277]=64483;
	multiplies[278]=64384;
	multiplies[279]=64280;
	multiplies[280]=64172;
	multiplies[281]=64060;
	multiplies[282]=63943;
	multiplies[283]=63821;
	multiplies[284]=63696;
	multiplies[285]=63566;
	multiplies[286]=63432;
	multiplies[287]=63293;
	multiplies[288]=63151;
	multiplies[289]=63004;
	multiplies[290]=62853;
	multiplies[291]=62698;
	multiplies[292]=62538;
	multiplies[293]=62375;
	multiplies[294]=62207;
	multiplies[295]=62036;
	multiplies[296]=61860;
	multiplies[297]=61680;
	multiplies[298]=61497;
	multiplies[299]=61309;
	multiplies[300]=61118;
	multiplies[301]=60922;
	multiplies[302]=60723;
	multiplies[303]=60519;
	multiplies[304]=60312;
	multiplies[305]=60102;
	multiplies[306]=59887;
	multiplies[307]=59669;
	multiplies[308]=59447;
	multiplies[309]=59221;
	multiplies[310]=58992;
	multiplies[311]=58759;
	multiplies[312]=58523;
	multiplies[313]=58283;
	multiplies[314]=58040;
	multiplies[315]=57793;
	multiplies[316]=57543;
	multiplies[317]=57289;
	multiplies[318]=57032;
	multiplies[319]=56772;
	multiplies[320]=56508;
	multiplies[321]=56242;
	multiplies[322]=55972;
	multiplies[323]=55699;
	multiplies[324]=55423;
	multiplies[325]=55144;
	multiplies[326]=54862;
	multiplies[327]=54577;
	multiplies[328]=54289;
	multiplies[329]=53998;
	multiplies[330]=53704;
	multiplies[331]=53408;
	multiplies[332]=53109;
	multiplies[333]=52807;
	multiplies[334]=52502;
	multiplies[335]=52195;
	multiplies[336]=51885;
	multiplies[337]=51573;
	multiplies[338]=51259;
	multiplies[339]=50941;
	multiplies[340]=50622;
	multiplies[341]=50300;
	multiplies[342]=49976;
	multiplies[343]=49650;
	multiplies[344]=49321;
	multiplies[345]=48991;
	multiplies[346]=48658;
	multiplies[347]=48324;
	multiplies[348]=47987;
	multiplies[349]=47648;
	multiplies[350]=47308;
	multiplies[351]=46966;
	multiplies[352]=46622;
	multiplies[353]=46276;
	multiplies[354]=45929;
	multiplies[355]=45580;
	multiplies[356]=45229;
	multiplies[357]=44877;
	multiplies[358]=44524;
	multiplies[359]=44169;
	multiplies[360]=43812;
	multiplies[361]=43455;
	multiplies[362]=43096;
	multiplies[363]=42736;
	multiplies[364]=42375;
	multiplies[365]=42013;
	multiplies[366]=41650;
	multiplies[367]=41286;
	multiplies[368]=40921;
	multiplies[369]=40555;
	multiplies[370]=40188;
	multiplies[371]=39821;
	multiplies[372]=39453;
	multiplies[373]=39084;
	multiplies[374]=38714;
	multiplies[375]=38345;
	multiplies[376]=37974;
	multiplies[377]=37604;
	multiplies[378]=37233;
	multiplies[379]=36861;
	multiplies[380]=36490;
	multiplies[381]=36118;
	multiplies[382]=35746;
	multiplies[383]=35374;
	multiplies[384]=35002;
	multiplies[385]=34630;
	multiplies[386]=34258;
	multiplies[387]=33886;
	multiplies[388]=33515;
	multiplies[389]=33144;
	multiplies[390]=32773;
	multiplies[391]=32402;
	multiplies[392]=32032;
	multiplies[393]=31663;
	multiplies[394]=31294;
	multiplies[395]=30925;
	multiplies[396]=30557;
	multiplies[397]=30190;
	multiplies[398]=29824;
	multiplies[399]=29459;
	multiplies[400]=29094;
	multiplies[401]=28730;
	multiplies[402]=28368;
	multiplies[403]=28006;
	multiplies[404]=27646;
	multiplies[405]=27286;
	multiplies[406]=26928;
	multiplies[407]=26571;
	multiplies[408]=26216;
	multiplies[409]=25861;
	multiplies[410]=25509;
	multiplies[411]=25157;
	multiplies[412]=24807;
	multiplies[413]=24459;
	multiplies[414]=24113;
	multiplies[415]=23768;
	multiplies[416]=23425;
	multiplies[417]=23083;
	multiplies[418]=22744;
	multiplies[419]=22406;
	multiplies[420]=22071;
	multiplies[421]=21737;
	multiplies[422]=21405;
	multiplies[423]=21076;
	multiplies[424]=20749;
	multiplies[425]=20423;
	multiplies[426]=20100;
	multiplies[427]=19780;
	multiplies[428]=19462;
	multiplies[429]=19146;
	multiplies[430]=18832;
	multiplies[431]=18521;
	multiplies[432]=18213;
	multiplies[433]=17907;
	multiplies[434]=17604;
	multiplies[435]=17303;
	multiplies[436]=17005;
	multiplies[437]=16710;
	multiplies[438]=16418;
	multiplies[439]=16129;
	multiplies[440]=15842;
	multiplies[441]=15559;
	multiplies[442]=15278;
	multiplies[443]=15000;
	multiplies[444]=14726;
	multiplies[445]=14455;
	multiplies[446]=14186;
	multiplies[447]=13921;
	multiplies[448]=13659;
	multiplies[449]=13401;
	multiplies[450]=13146;
	multiplies[451]=12894;
	multiplies[452]=12645;
	multiplies[453]=12400;
	multiplies[454]=12159;
	multiplies[455]=11920;
	multiplies[456]=11686;
	multiplies[457]=11455;
	multiplies[458]=11227;
	multiplies[459]=11004;
	multiplies[460]=10783;
	multiplies[461]=10567;
	multiplies[462]=10354;
	multiplies[463]=10145;
	multiplies[464]=9940;
	multiplies[465]=9739;
	multiplies[466]=9542;
	multiplies[467]=9348;
	multiplies[468]=9158;
	multiplies[469]=8973;
	multiplies[470]=8791;
	multiplies[471]=8613;
	multiplies[472]=8440;
	multiplies[473]=8270;
	multiplies[474]=8105;
	multiplies[475]=7943;
	multiplies[476]=7786;
	multiplies[477]=7633;
	multiplies[478]=7484;
	multiplies[479]=7339;
	multiplies[480]=7199;
	multiplies[481]=7062;
	multiplies[482]=6930;
	multiplies[483]=6803;
	multiplies[484]=6679;
	multiplies[485]=6560;
	multiplies[486]=6445;
	multiplies[487]=6335;
	multiplies[488]=6229;
	multiplies[489]=6128;
	multiplies[490]=6030;
	multiplies[491]=5938;
	multiplies[492]=5849;
	multiplies[493]=5765;
	multiplies[494]=5686;
	multiplies[495]=5611;
	multiplies[496]=5540;
	multiplies[497]=5474;
	multiplies[498]=5413;
	multiplies[499]=5356;
	multiplies[500]=5304;
	multiplies[501]=5256;
	multiplies[502]=5212;
	multiplies[503]=5174;
	multiplies[504]=5139;
	multiplies[505]=5110;
	multiplies[506]=5085;
	multiplies[507]=5064;
	multiplies[508]=5048;
	multiplies[509]=5036;
	multiplies[510]=5030;
	multiplies[511]=5027;

end



always@(posedge clk) 
	begin
		mul_out <= multiplies[mul_addr];
	end
	
endmodule
